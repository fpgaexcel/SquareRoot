program automatic test_program;
  import uvm_pkg::*;
endprogram
